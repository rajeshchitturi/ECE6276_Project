--Name of file : cordics.vhd

library ieee;